--asdf

-- another line