--asdf

